`timescale 1ns / 1ps
module SchoolSong(
    input beat,
	 input [1:0] func,
    input clk_5m,
    output reg [3:0] med = 4'b000,
    output reg[3:0] low = 4'b000
    );

reg [9:0] cnt;

always@(posedge beat )
begin
	 begin
	     if(cnt == 235 )
		      cnt <= 0;
		  else if(func[0] == 0 )
		      cnt <= 0;
			else
			cnt <= cnt + 1;
			case(cnt)
			0:{med,low} <= 'b0101_0000;    //��һ��
			1:{med,low} <= 'b0101_0000;
			2:{med,low} <= 'b0101_0000;
			3:{med,low} <= 'b0110_0000;
			
			4:{med,low} <= 'b0101_0000;
			5:{med,low} <= 'b0101_0000;
			6:{med,low} <= 'b0011_0000;
			7:{med,low} <= 'b0010_0000;
			
			8:{med,low} <= 'b0001_0000;
			9:{med,low} <= 'b0001_0000;
			10:{med,low} <= 'b0001_0000;
			11:{med,low} <= 'b0010_0000;
			
			12:{med,low} <= 'b0000_0101;
			13:{med,low} <= 'b0000_0101;
			14:{med,low} <= 'b0000_0000;
			15:{med,low} <= 'b0000_0101;
			
			16:{med,low} <= 'b0000_0110;
			17:{med,low} <= 'b0000_0110;
			18:{med,low} <= 'b0000_0101;
			19:{med,low} <= 'b0000_0101;
			
			20:{med,low} <= 'b0001_0000;
			21:{med,low} <= 'b0011_0000;
			22:{med,low} <= 'b0101_0000;
			23:{med,low} <= 'b0011_0000;
			
			24:{med,low} <= 'b0110_0000;
			25:{med,low} <= 'b0110_0000;
			26:{med,low} <= 'b0110_0000;
			27:{med,low} <= 'b0110_0000;
			
			28:{med,low} <= 'b0110_0000;
			29:{med,low} <= 'b0110_0000;
			30:{med,low} <= 'b0000_0000;
			31:{med,low} <= 'b0000_0000;
			
			32:{med,low} <= 'b0101_0000;  //�ڶ���
			33:{med,low} <= 'b0101_0000;
			34:{med,low} <= 'b0110_0000;
			35:{med,low} <= 'b0110_0000;
			
			36:{med,low} <= 'b0101_0000;
			37:{med,low} <= 'b0101_0000;
			38:{med,low} <= 'b0011_0000;
			39:{med,low} <= 'b0001_0000;
			
			40:{med,low} <= 'b0010_0000;
			41:{med,low} <= 'b0010_0000;
			42:{med,low} <= 'b0011_0000;
			43:{med,low} <= 'b0101_0000;
			
			44:{med,low} <= 'b0010_0000;
			45:{med,low} <= 'b0010_0000;
			46:{med,low} <= 'b0000_0000;
			47:{med,low} <= 'b0000_0000;
			
			48:{med,low} <= 'b0101_0000;
			49:{med,low} <= 'b0101_0000;
			50:{med,low} <= 'b0101_0000;
			51:{med,low} <= 'b0110_0000;
			
			52:{med,low} <= 'b0101_0000;
			53:{med,low} <= 'b0101_0000;
			54:{med,low} <= 'b0011_0000;
			55:{med,low} <= 'b0010_0000;
			
			56:{med,low} <= 'b0001_0000;
			57:{med,low} <= 'b0001_0000;
			58:{med,low} <= 'b0001_0000;
			59:{med,low} <= 'b0010_0000;
			
			60:{med,low} <= 'b0000_0101;
			61:{med,low} <= 'b0000_0101;
			62:{med,low} <= 'b0000_0000;
			63:{med,low} <= 'b0000_0000;
			
			64:{med,low} <= 'b0000_0110;    //������
			65:{med,low} <= 'b0000_0110;
			66:{med,low} <= 'b0000_0101;
			67:{med,low} <= 'b0000_0101;
			
			68:{med,low} <= 'b0001_0000;
			69:{med,low} <= 'b0011_0000;
			70:{med,low} <= 'b0101_0000;
			71:{med,low} <= 'b0110_0000;
			
			72:{med,low} <= 'b0011_0000;
			73:{med,low} <= 'b0011_0000;
			74:{med,low} <= 'b0011_0000;
			75:{med,low} <= 'b0011_0000;
			
			76:{med,low} <= 'b0011_0000;
			77:{med,low} <= 'b0011_0000;
			78:{med,low} <= 'b0000_0000;
			79:{med,low} <= 'b0000_0000;
			
			80:{med,low} <= 'b0101_0000;
			81:{med,low} <= 'b0101_0000;
			82:{med,low} <= 'b0101_0000;
			83:{med,low} <= 'b0110_0000;
			
			84:{med,low} <= 'b0101_0000;
			85:{med,low} <= 'b0101_0000;
			86:{med,low} <= 'b0101_0000;
			87:{med,low} <= 'b0011_0000;
			
			88:{med,low} <= 'b0010_0000;
			89:{med,low} <= 'b0010_0000;
			90:{med,low} <= 'b0011_0000;
			91:{med,low} <= 'b0110_0000;
			
			92:{med,low} <= 'b0101_0000;
			93:{med,low} <= 'b0101_0000;
			94:{med,low} <= 'b0000_0000;
			95:{med,low} <= 'b0000_0000;
			
			96:{med,low} <= 'b0011_0000;  //���ľ�
			97:{med,low} <= 'b0011_0000;
			98:{med,low} <= 'b0011_0000;
			99:{med,low} <= 'b0011_0000;
			
			100:{med,low} <= 'b0011_0000;
			101:{med,low} <= 'b0011_0000;
			102:{med,low} <= 'b0011_0000;
			103:{med,low} <= 'b0011_0000;
			
			104:{med,low} <= 'b0010_0000;
			105:{med,low} <= 'b0011_0000;
			106:{med,low} <= 'b0010_0000;
			107:{med,low} <= 'b0001_0000;
			
			108:{med,low} <= 'b0000_0110;
			109:{med,low} <= 'b0000_0110;
			110:{med,low} <= 'b0000_0000;
			111:{med,low} <= 'b0000_0101;
			
			112:{med,low} <= 'b0001_0000;
			113:{med,low} <= 'b0011_0000;
			114:{med,low} <= 'b0101_0000;
			115:{med,low} <= 'b0110_0000;
			
			116:{med,low} <= 'b0101_0000;
			117:{med,low} <= 'b0101_0000;
			118:{med,low} <= 'b0000_0000;
			119:{med,low} <= 'b0000_0000;
			
			120:{med,low} <= 'b0010_0000;
			121:{med,low} <= 'b0011_0000;
			122:{med,low} <= 'b0010_0000;
			123:{med,low} <= 'b0001_0000;
			
			124:{med,low} <= 'b0010_0000;
			125:{med,low} <= 'b0010_0000;
			126:{med,low} <= 'b0000_0000;
			127:{med,low} <= 'b0000_0101;
			
			128:{med,low} <= 'b0011_0000;    //�����
			129:{med,low} <= 'b0011_0000;
			130:{med,low} <= 'b0011_0000;
			131:{med,low} <= 'b0011_0000;
			
			132:{med,low} <= 'b0010_0000;
			133:{med,low} <= 'b0010_0000;
			134:{med,low} <= 'b0011_0000;
			135:{med,low} <= 'b0011_0000;
			
			136:{med,low} <= 'b0010_0000;
			137:{med,low} <= 'b0011_0000;
			138:{med,low} <= 'b0010_0000;
			139:{med,low} <= 'b0001_0000;
			
			140:{med,low} <= 'b0000_0110;
			141:{med,low} <= 'b0000_0110;
			142:{med,low} <= 'b0000_0000;
			143:{med,low} <= 'b0000_0101;
			
			144:{med,low} <= 'b0101_0000;
			145:{med,low} <= 'b0101_0000;
			146:{med,low} <= 'b0101_0000;
			147:{med,low} <= 'b0101_0000;
			
			148:{med,low} <= 'b0110_0000;
			149:{med,low} <= 'b0110_0000;
			150:{med,low} <= 'b0110_0000;
			151:{med,low} <= 'b0110_0000;
			
			152:{med,low} <= 'b0101_0000;
			153:{med,low} <= 'b0101_0000;
			154:{med,low} <= 'b0010_0000;
			155:{med,low} <= 'b0010_0000;
			
			156:{med,low} <= 'b0101_0000;
			157:{med,low} <= 'b0101_0000;
			158:{med,low} <= 'b0101_0000;
			159:{med,low} <= 'b0101_0000;
			
			160:{med,low} <= 'b0110_0000;   //������
			161:{med,low} <= 'b0110_0000;
			162:{med,low} <= 'b0101_0000;
			163:{med,low} <= 'b0110_0000;
			
			164:{med,low} <= 'b0011_0000;
			165:{med,low} <= 'b0011_0000;
			166:{med,low} <= 'b0000_0000;
			167:{med,low} <= 'b0000_0000;
			
			168:{med,low} <= 'b0010_0000;
			169:{med,low} <= 'b0101_0000;
			170:{med,low} <= 'b0011_0000;
			171:{med,low} <= 'b0001_0000;
			
			172:{med,low} <= 'b0010_0000;
			173:{med,low} <= 'b0010_0000;
			174:{med,low} <= 'b0000_0000;
			175:{med,low} <= 'b0000_0000;
			
			176:{med,low} <= 'b0000_0101;
			177:{med,low} <= 'b0000_0000;
			178:{med,low} <= 'b0001_0000;
			179:{med,low} <= 'b0000_0000;
			
			180:{med,low} <= 'b0101_0000;
			181:{med,low} <= 'b0000_0000;
			182:{med,low} <= 'b0011_0000;
			183:{med,low} <= 'b0000_0000;
			
			184:{med,low} <= 'b0010_0000;
			185:{med,low} <= 'b0010_0000;
			186:{med,low} <= 'b0110_0000;
			187:{med,low} <= 'b0110_0000;
			
			188:{med,low} <= 'b0101_0000;
			189:{med,low} <= 'b0101_0000;
			190:{med,low} <= 'b0000_0000;
			191:{med,low} <= 'b0000_0000;
			
			192:{med,low} <= 'b0110_0000;    //���߾�
			193:{med,low} <= 'b0110_0000;
			194:{med,low} <= 'b0110_0000;
			195:{med,low} <= 'b0110_0000;
			
			196:{med,low} <= 'b0101_0000;
			197:{med,low} <= 'b0101_0000;
			198:{med,low} <= 'b0110_0000;
			199:{med,low} <= 'b0110_0000;
			
			200:{med,low} <= 'b0101_0000;
			201:{med,low} <= 'b0101_0000;
			202:{med,low} <= 'b0011_0000;
			203:{med,low} <= 'b0001_0000;
			
			204:{med,low} <= 'b0010_0000;
			205:{med,low} <= 'b0010_0000;
			206:{med,low} <= 'b0000_0110;
			207:{med,low} <= 'b0000_0101;
			
			208:{med,low} <= 'b0001_0000;
			209:{med,low} <= 'b0000_0000;
			210:{med,low} <= 'b0010_0000;
			211:{med,low} <= 'b0000_0000;
			
			212:{med,low} <= 'b0011_0000;
			213:{med,low} <= 'b0000_0000;
			214:{med,low} <= 'b0101_0000;
			215:{med,low} <= 'b0000_0000;
			
			216:{med,low} <= 'b0110_0000;
			217:{med,low} <= 'b0110_0000;
			218:{med,low} <= 'b0110_0000;
			219:{med,low} <= 'b0110_0000;
			
			220:{med,low} <= 'b0101_0000;
			221:{med,low} <= 'b0101_0000;
			222:{med,low} <= 'b0101_0000;
			223:{med,low} <= 'b0101_0000;
			
			224:{med,low} <= 'b0101_0000;
			225:{med,low} <= 'b0101_0000;
			226:{med,low} <= 'b0101_0000;
			227:{med,low} <= 'b0101_0000;
			
			228:{med,low} <= 'b0000_0000;
			229:{med,low} <= 'b0000_0000;
			230:{med,low} <= 'b0000_0000;
			231:{med,low} <= 'b0000_0000;
			
			232:{med,low} <= 'b0000_0000;
			233:{med,low} <= 'b0000_0000;
			234:{med,low} <= 'b0000_0000;
			235:{med,low} <= 'b0000_0000;
			endcase
	 end
end

endmodule
