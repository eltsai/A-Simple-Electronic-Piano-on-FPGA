`timescale 1ns / 1ps
module WaterLight(       //��ˮ��ģ��
    input           beat,
    input     [3:0] func,
    output reg[7:0] L,
    input           rst_n
    );
	 
reg [7:0] cnt = 0;	 
	 
always@(posedge beat)
begin
    if(~rst_n)
	 L <= 8'b0;
	 else if(func == 2'b11)
	 L <= 8'b0;
	 else if(func == 2'b00)
	 L <= 8'b0; 
	 else
	 begin
	     case(cnt)
	     0: L <= 8'b0000_0001;
	     1: L <= 8'b0000_0010;
    	  2: L <= 8'b0000_0100;
	     3: L <= 8'b0000_1000;
	     4: L <= 8'b0001_0000;
	     5: L <= 8'b0010_0000;
	     6: L <= 8'b0100_0000;
	     7: L <= 8'b1000_0000;
		  
		  8: L <= 8'b1000_0000;
		  9: L <= 8'b0100_0000;
		  10: L <= 8'b0010_0000;
		  11: L <= 8'b0001_0000;
		  12: L <= 8'b0000_1000;
		  13: L <= 8'b0000_0100;
		  14: L <= 8'b0000_0010;
		  15: L <= 8'b0000_0001;
		  
		  16: L <= 8'b0001_1000;
        17: L <= 8'b0010_0100;
        18: L <= 8'b0100_0010;
        19: L <= 8'b1000_0001;
        20: L <= 8'b1000_0001;
        21: L <= 8'b0100_0010;
        22: L <= 8'b0010_0100;
        23: L <= 8'b0001_1000; 

		  24: L <= 8'b0001_1000;
        25: L <= 8'b0010_0100;
        26: L <= 8'b0100_0010;
        27: L <= 8'b1000_0001;
        28: L <= 8'b1000_0001;
        29: L <= 8'b0100_0010;
        30: L <= 8'b0010_0100;
        31: L <= 8'b0001_1000; 		  
	    
		 default: L <= 8'b0000_0000;
	 endcase
	 if(cnt == 8'h31)
	     cnt <= 0;
	 else 
	     cnt <= cnt + 1;
	 end
	 

end

endmodule
